
`timescale 1ps/1ps
module bm_ce_rom (clock, addr, rdata);

input              clock    ;
input  [7:0]       addr     ;
output [64:0]      rdata    ;

reg    [64:0]      rdata    ;

always @(posedge clock)
  case(addr)
    8'd0: rdata <= #1 {30'd1, 22'd4194292, 13'd8160};
    8'd1: rdata <= #1 {30'd4186134, 22'd4177972, 13'd8097};
    8'd2: rdata <= #1 {30'd8356010, 22'd4161778, 13'd8034};
    8'd3: rdata <= #1 {30'd12509756, 22'd4145710, 13'd7973};
    8'd4: rdata <= #1 {30'd16647494, 22'd4129765, 13'd7911};
    8'd5: rdata <= #1 {30'd20769349, 22'd4113942, 13'd7851};
    8'd6: rdata <= #1 {30'd24875441, 22'd4098240, 13'd7791};
    8'd7: rdata <= #1 {30'd28965891, 22'd4082658, 13'd7732};
    8'd8: rdata <= #1 {30'd33040818, 22'd4067193, 13'd7674};
    8'd9: rdata <= #1 {30'd37100338, 22'd4051845, 13'd7616};
    8'd10: rdata <= #1 {30'd41144568, 22'd4036613, 13'd7559};
    8'd11: rdata <= #1 {30'd45173623, 22'd4021494, 13'd7503};
    8'd12: rdata <= #1 {30'd49187615, 22'd4006489, 13'd7447};
    8'd13: rdata <= #1 {30'd53186658, 22'd3991595, 13'd7392};
    8'd14: rdata <= #1 {30'd57170863, 22'd3976811, 13'd7337};
    8'd15: rdata <= #1 {30'd61140338, 22'd3962137, 13'd7283};
    8'd16: rdata <= #1 {30'd65095193, 22'd3947570, 13'd7230};
    8'd17: rdata <= #1 {30'd69035534, 22'd3933110, 13'd7177};
    8'd18: rdata <= #1 {30'd72961468, 22'd3918756, 13'd7125};
    8'd19: rdata <= #1 {30'd76873100, 22'd3904506, 13'd7073};
    8'd20: rdata <= #1 {30'd80770534, 22'd3890359, 13'd7022};
    8'd21: rdata <= #1 {30'd84653872, 22'd3876315, 13'd6972};
    8'd22: rdata <= #1 {30'd88523216, 22'd3862371, 13'd6922};
    8'd23: rdata <= #1 {30'd92378667, 22'd3848528, 13'd6872};
    8'd24: rdata <= #1 {30'd96220323, 22'd3834783, 13'd6823};
    8'd25: rdata <= #1 {30'd100048284, 22'd3821136, 13'd6775};
    8'd26: rdata <= #1 {30'd103862646, 22'd3807586, 13'd6727};
    8'd27: rdata <= #1 {30'd107663506, 22'd3794132, 13'd6680};
    8'd28: rdata <= #1 {30'd111450959, 22'd3780772, 13'd6633};
    8'd29: rdata <= #1 {30'd115225099, 22'd3767507, 13'd6587};
    8'd30: rdata <= #1 {30'd118986020, 22'd3754333, 13'd6541};
    8'd31: rdata <= #1 {30'd122733814, 22'd3741252, 13'd6495};
    8'd32: rdata <= #1 {30'd126468572, 22'd3728262, 13'd6450};
    8'd33: rdata <= #1 {30'd130190384, 22'd3715361, 13'd6406};
    8'd34: rdata <= #1 {30'd133899341, 22'd3702550, 13'd6362};
    8'd35: rdata <= #1 {30'd137595530, 22'd3689826, 13'd6318};
    8'd36: rdata <= #1 {30'd141279039, 22'd3677190, 13'd6275};
    8'd37: rdata <= #1 {30'd144949955, 22'd3664640, 13'd6232};
    8'd38: rdata <= #1 {30'd148608363, 22'd3652175, 13'd6190};
    8'd39: rdata <= #1 {30'd152254349, 22'd3639795, 13'd6148};
    8'd40: rdata <= #1 {30'd155887997, 22'd3627498, 13'd6107};
    8'd41: rdata <= #1 {30'd159509389, 22'd3615285, 13'd6066};
    8'd42: rdata <= #1 {30'd163118608, 22'd3603153, 13'd6025};
    8'd43: rdata <= #1 {30'd166715737, 22'd3591102, 13'd5985};
    8'd44: rdata <= #1 {30'd170300855, 22'd3579132, 13'd5945};
    8'd45: rdata <= #1 {30'd173874042, 22'd3567241, 13'd5906};
    8'd46: rdata <= #1 {30'd177435378, 22'd3555429, 13'd5867};
    8'd47: rdata <= #1 {30'd180984941, 22'd3543695, 13'd5828};
    8'd48: rdata <= #1 {30'd184522809, 22'd3532038, 13'd5790};
    8'd49: rdata <= #1 {30'd188049058, 22'd3520458, 13'd5752};
    8'd50: rdata <= #1 {30'd191563764, 22'd3508953, 13'd5715};
    8'd51: rdata <= #1 {30'd195067003, 22'd3497523, 13'd5678};
    8'd52: rdata <= #1 {30'd198558849, 22'd3486168, 13'd5641};
    8'd53: rdata <= #1 {30'd202039377, 22'd3474886, 13'd5605};
    8'd54: rdata <= #1 {30'd205508659, 22'd3463677, 13'd5569};
    8'd55: rdata <= #1 {30'd208966768, 22'd3452539, 13'd5533};
    8'd56: rdata <= #1 {30'd212413775, 22'd3441474, 13'd5498};
    8'd57: rdata <= #1 {30'd215849752, 22'd3430479, 13'd5463};
    8'd58: rdata <= #1 {30'd219274768, 22'd3419553, 13'd5428};
    8'd59: rdata <= #1 {30'd222688895, 22'd3408698, 13'd5394};
    8'd60: rdata <= #1 {30'd226092200, 22'd3397911, 13'd5359};
    8'd61: rdata <= #1 {30'd229484752, 22'd3387192, 13'd5326};
    8'd62: rdata <= #1 {30'd232866618, 22'd3376540, 13'd5292};
    8'd63: rdata <= #1 {30'd236237867, 22'd3365956, 13'd5259};
    8'd64: rdata <= #1 {30'd239598564, 22'd3355437, 13'd5227};
    8'd65: rdata <= #1 {30'd242948775, 22'd3344984, 13'd5194};
    8'd66: rdata <= #1 {30'd246288566, 22'd3334596, 13'd5162};
    8'd67: rdata <= #1 {30'd249618001, 22'd3324272, 13'd5130};
    8'd68: rdata <= #1 {30'd252937143, 22'd3314012, 13'd5098};
    8'd69: rdata <= #1 {30'd256246058, 22'd3303815, 13'd5067};
    8'd70: rdata <= #1 {30'd259544806, 22'd3293681, 13'd5036};
    8'd71: rdata <= #1 {30'd262833451, 22'd3283608, 13'd5006};
    8'd72: rdata <= #1 {30'd266112055, 22'd3273597, 13'd4975};
    8'd73: rdata <= #1 {30'd269380678, 22'd3263647, 13'd4945};
    8'd74: rdata <= #1 {30'd272639381, 22'd3253758, 13'd4915};
    8'd75: rdata <= #1 {30'd275888224, 22'd3243927, 13'd4885};
    8'd76: rdata <= #1 {30'd279127267, 22'd3234157, 13'd4856};
    8'd77: rdata <= #1 {30'd282356568, 22'd3224444, 13'd4827};
    8'd78: rdata <= #1 {30'd285576186, 22'd3214790, 13'd4798};
    8'd79: rdata <= #1 {30'd288786179, 22'd3205194, 13'd4770};
    8'd80: rdata <= #1 {30'd291986604, 22'd3195655, 13'd4741};
    8'd81: rdata <= #1 {30'd295177518, 22'd3186172, 13'd4713};
    8'd82: rdata <= #1 {30'd298358978, 22'd3176746, 13'd4685};
    8'd83: rdata <= #1 {30'd301531039, 22'd3167375, 13'd4658};
    8'd84: rdata <= #1 {30'd304693756, 22'd3158059, 13'd4631};
    8'd85: rdata <= #1 {30'd307847185, 22'd3148798, 13'd4604};
    8'd86: rdata <= #1 {30'd310991380, 22'd3139591, 13'd4577};
    8'd87: rdata <= #1 {30'd314126395, 22'd3130438, 13'd4550};
    8'd88: rdata <= #1 {30'd317252283, 22'd3121338, 13'd4524};
    8'd89: rdata <= #1 {30'd320369098, 22'd3112290, 13'd4498};
    8'd90: rdata <= #1 {30'd323476891, 22'd3103295, 13'd4472};
    8'd91: rdata <= #1 {30'd326575715, 22'd3094352, 13'd4446};
    8'd92: rdata <= #1 {30'd329665622, 22'd3085460, 13'd4420};
    8'd93: rdata <= #1 {30'd332746662, 22'd3076619, 13'd4395};
    8'd94: rdata <= #1 {30'd335818887, 22'd3067829, 13'd4370};
    8'd95: rdata <= #1 {30'd338882346, 22'd3059089, 13'd4345};
    8'd96: rdata <= #1 {30'd341937090, 22'd3050398, 13'd4321};
    8'd97: rdata <= #1 {30'd344983168, 22'd3041757, 13'd4296};
    8'd98: rdata <= #1 {30'd348020630, 22'd3033164, 13'd4272};
    8'd99: rdata <= #1 {30'd351049523, 22'd3024620, 13'd4248};
    8'd100: rdata <= #1 {30'd354069895, 22'd3016124, 13'd4224};
    8'd101: rdata <= #1 {30'd357081796, 22'd3007676, 13'd4201};
    8'd102: rdata <= #1 {30'd360085271, 22'd2999274, 13'd4177};
    8'd103: rdata <= #1 {30'd363080369, 22'd2990920, 13'd4154};
    8'd104: rdata <= #1 {30'd366067136, 22'd2982612, 13'd4131};
    8'd105: rdata <= #1 {30'd369045617, 22'd2974350, 13'd4108};
    8'd106: rdata <= #1 {30'd372015859, 22'd2966133, 13'd4086};
    8'd107: rdata <= #1 {30'd374977907, 22'd2957962, 13'd4063};
    8'd108: rdata <= #1 {30'd377931807, 22'd2949836, 13'd4041};
    8'd109: rdata <= #1 {30'd380877602, 22'd2941754, 13'd4019};
    8'd110: rdata <= #1 {30'd383815338, 22'd2933717, 13'd3997};
    8'd111: rdata <= #1 {30'd386745059, 22'd2925723, 13'd3975};
    8'd112: rdata <= #1 {30'd389666807, 22'd2917773, 13'd3954};
    8'd113: rdata <= #1 {30'd392580626, 22'd2909865, 13'd3932};
    8'd114: rdata <= #1 {30'd395486560, 22'd2902001, 13'd3911};
    8'd115: rdata <= #1 {30'd398384650, 22'd2894179, 13'd3890};
    8'd116: rdata <= #1 {30'd401274940, 22'd2886399, 13'd3869};
    8'd117: rdata <= #1 {30'd404157470, 22'd2878661, 13'd3848};
    8'd118: rdata <= #1 {30'd407032282, 22'd2870964, 13'd3828};
    8'd119: rdata <= #1 {30'd409899418, 22'd2863308, 13'd3808};
    8'd120: rdata <= #1 {30'd412758919, 22'd2855693, 13'd3787};
    8'd121: rdata <= #1 {30'd415610825, 22'd2848118, 13'd3767};
    8'd122: rdata <= #1 {30'd418455175, 22'd2840583, 13'd3747};
    8'd123: rdata <= #1 {30'd421292011, 22'd2833088, 13'd3728};
    8'd124: rdata <= #1 {30'd424121372, 22'd2825633, 13'd3708};
    8'd125: rdata <= #1 {30'd426943297, 22'd2818216, 13'd3689};
    8'd126: rdata <= #1 {30'd429757825, 22'd2810839, 13'd3670};
    8'd127: rdata <= #1 {30'd432564995, 22'd2803500, 13'd3650};
    8'd128: rdata <= #1 {30'd435364845, 22'd2796199, 13'd3631};
    8'd129: rdata <= #1 {30'd438157413, 22'd2788936, 13'd3613};
    8'd130: rdata <= #1 {30'd440942737, 22'd2781711, 13'd3594};
    8'd131: rdata <= #1 {30'd443720855, 22'd2774523, 13'd3575};
    8'd132: rdata <= #1 {30'd446491803, 22'd2767372, 13'd3557};
    8'd133: rdata <= #1 {30'd449255619, 22'd2760258, 13'd3539};
    8'd134: rdata <= #1 {30'd452012339, 22'd2753181, 13'd3521};
    8'd135: rdata <= #1 {30'd454761999, 22'd2746139, 13'd3503};
    8'd136: rdata <= #1 {30'd457504636, 22'd2739134, 13'd3485};
    8'd137: rdata <= #1 {30'd460240285, 22'd2732164, 13'd3467};
    8'd138: rdata <= #1 {30'd462968983, 22'd2725230, 13'd3450};
    8'd139: rdata <= #1 {30'd465690763, 22'd2718330, 13'd3432};
    8'd140: rdata <= #1 {30'd468405662, 22'd2711466, 13'd3415};
    8'd141: rdata <= #1 {30'd471113713, 22'd2704636, 13'd3398};
    8'd142: rdata <= #1 {30'd473814952, 22'd2697841, 13'd3381};
    8'd143: rdata <= #1 {30'd476509412, 22'd2691079, 13'd3364};
    8'd144: rdata <= #1 {30'd479197128, 22'd2684351, 13'd3347};
    8'd145: rdata <= #1 {30'd481878132, 22'd2677657, 13'd3330};
    8'd146: rdata <= #1 {30'd484552460, 22'd2670996, 13'd3314};
    8'd147: rdata <= #1 {30'd487220143, 22'd2664369, 13'd3297};
    8'd148: rdata <= #1 {30'd489881214, 22'd2657774, 13'd3281};
    8'd149: rdata <= #1 {30'd492535707, 22'd2651211, 13'd3265};
    8'd150: rdata <= #1 {30'd495183654, 22'd2644681, 13'd3249};
    8'd151: rdata <= #1 {30'd497825086, 22'd2638183, 13'd3233};
    8'd152: rdata <= #1 {30'd500460037, 22'd2631717, 13'd3217};
    8'd153: rdata <= #1 {30'd503088537, 22'd2625283, 13'd3202};
    8'd154: rdata <= #1 {30'd505710619, 22'd2618880, 13'd3186};
    8'd155: rdata <= #1 {30'd508326312, 22'd2612508, 13'd3171};
    8'd156: rdata <= #1 {30'd510935650, 22'd2606167, 13'd3155};
    8'd157: rdata <= #1 {30'd513538662, 22'd2599856, 13'd3140};
    8'd158: rdata <= #1 {30'd516135378, 22'd2593576, 13'd3125};
    8'd159: rdata <= #1 {30'd518725830, 22'd2587327, 13'd3110};
    8'd160: rdata <= #1 {30'd521310048, 22'd2581107, 13'd3095};
    8'd161: rdata <= #1 {30'd523888061, 22'd2574918, 13'd3080};
    8'd162: rdata <= #1 {30'd526459899, 22'd2568758, 13'd3065};
    8'd163: rdata <= #1 {30'd529025591, 22'd2562627, 13'd3051};
    8'd164: rdata <= #1 {30'd531585167, 22'd2556525, 13'd3036};
    8'd165: rdata <= #1 {30'd534138657, 22'd2550453, 13'd3022};
    8'd166: rdata <= #1 {30'd536686088, 22'd2544409, 13'd3008};
    8'd167: rdata <= #1 {30'd539227491, 22'd2538394, 13'd2993};
    8'd168: rdata <= #1 {30'd541762892, 22'd2532407, 13'd2979};
    8'd169: rdata <= #1 {30'd544292320, 22'd2526449, 13'd2965};
    8'd170: rdata <= #1 {30'd546815804, 22'd2520518, 13'd2951};
    8'd171: rdata <= #1 {30'd549333370, 22'd2514615, 13'd2938};
    8'd172: rdata <= #1 {30'd551845048, 22'd2508740, 13'd2924};
    8'd173: rdata <= #1 {30'd554350865, 22'd2502892, 13'd2910};
    8'd174: rdata <= #1 {30'd556850847, 22'd2497071, 13'd2897};
    8'd175: rdata <= #1 {30'd559345022, 22'd2491278, 13'd2883};
    8'd176: rdata <= #1 {30'd561833416, 22'd2485511, 13'd2870};
    8'd177: rdata <= #1 {30'd564316058, 22'd2479771, 13'd2857};
    8'd178: rdata <= #1 {30'd566792972, 22'd2474057, 13'd2844};
    8'd179: rdata <= #1 {30'd569264185, 22'd2468370, 13'd2831};
    8'd180: rdata <= #1 {30'd571729724, 22'd2462708, 13'd2818};
    8'd181: rdata <= #1 {30'd574189615, 22'd2457073, 13'd2805};
    8'd182: rdata <= #1 {30'd576643883, 22'd2451463, 13'd2792};
    8'd183: rdata <= #1 {30'd579092555, 22'd2445879, 13'd2779};
    8'd184: rdata <= #1 {30'd581535654, 22'd2440320, 13'd2767};
    8'd185: rdata <= #1 {30'd583973207, 22'd2434786, 13'd2754};
    8'd186: rdata <= #1 {30'd586405240, 22'd2429278, 13'd2742};
    8'd187: rdata <= #1 {30'd588831776, 22'd2423794, 13'd2729};
    8'd188: rdata <= #1 {30'd591252841, 22'd2418335, 13'd2717};
    8'd189: rdata <= #1 {30'd593668459, 22'd2412901, 13'd2705};
    8'd190: rdata <= #1 {30'd596078655, 22'd2407491, 13'd2693};
    8'd191: rdata <= #1 {30'd598483453, 22'd2402105, 13'd2681};
    8'd192: rdata <= #1 {30'd600882877, 22'd2396743, 13'd2669};
    8'd193: rdata <= #1 {30'd603276951, 22'd2391405, 13'd2657};
    8'd194: rdata <= #1 {30'd605665699, 22'd2386091, 13'd2645};
    8'd195: rdata <= #1 {30'd608049145, 22'd2380800, 13'd2634};
    8'd196: rdata <= #1 {30'd610427312, 22'd2375533, 13'd2622};
    8'd197: rdata <= #1 {30'd612800223, 22'd2370289, 13'd2610};
    8'd198: rdata <= #1 {30'd615167901, 22'd2365068, 13'd2599};
    8'd199: rdata <= #1 {30'd617530370, 22'd2359870, 13'd2588};
    8'd200: rdata <= #1 {30'd619887653, 22'd2354695, 13'd2576};
    8'd201: rdata <= #1 {30'd622239772, 22'd2349542, 13'd2565};
    8'd202: rdata <= #1 {30'd624586750, 22'd2344412, 13'd2554};
    8'd203: rdata <= #1 {30'd626928609, 22'd2339305, 13'd2543};
    8'd204: rdata <= #1 {30'd629265371, 22'd2334219, 13'd2532};
    8'd205: rdata <= #1 {30'd631597058, 22'd2329156, 13'd2521};
    8'd206: rdata <= #1 {30'd633923694, 22'd2324114, 13'd2510};
    8'd207: rdata <= #1 {30'd636245299, 22'd2319095, 13'd2499};
    8'd208: rdata <= #1 {30'd638561895, 22'd2314097, 13'd2488};
    8'd209: rdata <= #1 {30'd640873503, 22'd2309120, 13'd2478};
    8'd210: rdata <= #1 {30'd643180146, 22'd2304165, 13'd2467};
    8'd211: rdata <= #1 {30'd645481844, 22'd2299231, 13'd2456};
    8'd212: rdata <= #1 {30'd647778619, 22'd2294318, 13'd2446};
    8'd213: rdata <= #1 {30'd650070492, 22'd2289426, 13'd2436};
    8'd214: rdata <= #1 {30'd652357482, 22'd2284555, 13'd2425};
    8'd215: rdata <= #1 {30'd654639613, 22'd2279705, 13'd2415};
    8'd216: rdata <= #1 {30'd656916903, 22'd2274875, 13'd2405};
    8'd217: rdata <= #1 {30'd659189373, 22'd2270065, 13'd2395};
    8'd218: rdata <= #1 {30'd661457044, 22'd2265276, 13'd2385};
    8'd219: rdata <= #1 {30'd663719936, 22'd2260507, 13'd2374};
    8'd220: rdata <= #1 {30'd665978069, 22'd2255758, 13'd2365};
    8'd221: rdata <= #1 {30'd668231463, 22'd2251029, 13'd2355};
    8'd222: rdata <= #1 {30'd670480138, 22'd2246320, 13'd2345};
    8'd223: rdata <= #1 {30'd672724113, 22'd2241630, 13'd2335};
    8'd224: rdata <= #1 {30'd674963409, 22'd2236960, 13'd2325};
    8'd225: rdata <= #1 {30'd677198044, 22'd2232310, 13'd2316};
    8'd226: rdata <= #1 {30'd679428038, 22'd2227678, 13'd2306};
    8'd227: rdata <= #1 {30'd681653411, 22'd2223066, 13'd2297};
    8'd228: rdata <= #1 {30'd683874180, 22'd2218473, 13'd2287};
    8'd229: rdata <= #1 {30'd686090367, 22'd2213899, 13'd2278};
    8'd230: rdata <= #1 {30'd688301988, 22'd2209344, 13'd2268};
    8'd231: rdata <= #1 {30'd690509063, 22'd2204807, 13'd2259};
    8'd232: rdata <= #1 {30'd692711611, 22'd2200289, 13'd2250};
    8'd233: rdata <= #1 {30'd694909651, 22'd2195789, 13'd2241};
    8'd234: rdata <= #1 {30'd697103200, 22'd2191308, 13'd2231};
    8'd235: rdata <= #1 {30'd699292277, 22'd2186845, 13'd2222};
    8'd236: rdata <= #1 {30'd701476900, 22'd2182400, 13'd2213};
    8'd237: rdata <= #1 {30'd703657087, 22'd2177974, 13'd2204};
    8'd238: rdata <= #1 {30'd705832856, 22'd2173565, 13'd2196};
    8'd239: rdata <= #1 {30'd708004225, 22'd2169174, 13'd2187};
    8'd240: rdata <= #1 {30'd710171213, 22'd2164800, 13'd2178};
    8'd241: rdata <= #1 {30'd712333836, 22'd2160445, 13'd2169};
    8'd242: rdata <= #1 {30'd714492111, 22'd2156106, 13'd2160};
    8'd243: rdata <= #1 {30'd716646057, 22'd2151786, 13'd2152};
    8'd244: rdata <= #1 {30'd718795691, 22'd2147482, 13'd2143};
    8'd245: rdata <= #1 {30'd720941031, 22'd2143196, 13'd2135};
    8'd246: rdata <= #1 {30'd723082092, 22'd2138926, 13'd2126};
    8'd247: rdata <= #1 {30'd725218892, 22'd2134674, 13'd2118};
    8'd248: rdata <= #1 {30'd727351449, 22'd2130439, 13'd2109};
    8'd249: rdata <= #1 {30'd729479778, 22'd2126220, 13'd2101};
    8'd250: rdata <= #1 {30'd731603897, 22'd2122018, 13'd2093};
    8'd251: rdata <= #1 {30'd733723822, 22'd2117832, 13'd2084};
    8'd252: rdata <= #1 {30'd735839570, 22'd2113663, 13'd2076};
    8'd253: rdata <= #1 {30'd737951158, 22'd2109511, 13'd2068};
    8'd254: rdata <= #1 {30'd740058601, 22'd2105375, 13'd2060};
    8'd255: rdata <= #1 {30'd742161915, 22'd2101255, 13'd2052};
    default: rdata <= #1 65'd0;
  endcase

endmodule

